library verilog;
use verilog.vl_types.all;
entity tb_MBE_encoder is
end tb_MBE_encoder;
