library verilog;
use verilog.vl_types.all;
entity tb_RISC is
end tb_RISC;
