LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY instruction_memory IS
PORT(
		CLK, MEM_READ: IN STD_LOGIC;
		ADDR: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_OUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END instruction_memory;

ARCHITECTURE structure OF instruction_memory IS

type MEM_TYP IS ARRAY(4194300 TO 4194428) OF STD_LOGIC_VECTOR(7 DOWNTO 0); --LARGER MEMORY TO STORE THE NOP
SIGNAL IM: MEM_TYP;
--SIGNAL DATA_OUT_s: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

IM(4194304) <= "00010011";
IM(4194305) <= "00001000";
IM(4194306) <= "01110000";
IM(4194307) <= "00000000";
IM(4194308) <= "00010111";
IM(4194309) <= "00000010";
IM(4194310) <= "11000001";
IM(4194311) <= "00001111";
IM(4194312) <= "00010011";
IM(4194313) <= "00000010";
IM(4194314) <= "11000010";
IM(4194315) <= "11111111";
IM(4194316) <= "10010111";
IM(4194317) <= "00000010";
IM(4194318) <= "11000001";
IM(4194319) <= "00001111";
IM(4194320) <= "10010011";
IM(4194321) <= "10000010";
IM(4194322) <= "00000010";
IM(4194323) <= "00000001";
IM(4194324) <= "10110111";
IM(4194325) <= "00000110";
IM(4194326) <= "00000000";
IM(4194327) <= "01000000";
IM(4194328) <= "10010011";
IM(4194329) <= "10000110";
IM(4194330) <= "11110110";
IM(4194331) <= "11111111";
IM(4194332) <= "01100011";
IM(4194333) <= "00000110";
IM(4194334) <= "00001000";
IM(4194335) <= "00000100";
IM(4194336) <= "00000011";
IM(4194337) <= "00100100";
IM(4194338) <= "00000010";
IM(4194339) <= "00000000";
IM(4194340) <= "00010011";
IM(4194341) <= "00000000";
IM(4194342) <= "00000000";
IM(4194343) <= "00000000";
IM(4194344) <= "10010011";
IM(4194345) <= "01010100";
IM(4194346) <= "11110100";
IM(4194347) <= "01000001";
IM(4194348) <= "00110011";
IM(4194349) <= "01000101";
IM(4194350) <= "10010100";
IM(4194351) <= "00000000";
IM(4194352) <= "10010011";
IM(4194353) <= "11110100";
IM(4194354) <= "00010100";
IM(4194355) <= "00000000";
IM(4194356) <= "00110011";
IM(4194357) <= "00000101";
IM(4194358) <= "10010101";
IM(4194359) <= "00000000";
IM(4194360) <= "00010011";
IM(4194361) <= "00000010";
IM(4194362) <= "01000010";
IM(4194363) <= "00000000";
IM(4194364) <= "00010011";
IM(4194365) <= "00001000";
IM(4194366) <= "11111000";
IM(4194367) <= "11111111";
IM(4194368) <= "10110011";
IM(4194369) <= "00100101";
IM(4194370) <= "11010101";
IM(4194371) <= "00000000";
IM(4194372) <= "11100011";
IM(4194373) <= "10001100";
IM(4194374) <= "00000101";
IM(4194375) <= "11111100";
IM(4194376) <= "00010011";
IM(4194377) <= "00000000";
IM(4194378) <= "00000000";
IM(4194379) <= "00000000";
IM(4194380) <= "00010011";
IM(4194381) <= "00000000";
IM(4194382) <= "00000000";
IM(4194383) <= "00000000";
IM(4194384) <= "00010011";
IM(4194385) <= "00000000";
IM(4194386) <= "00000000";
IM(4194387) <= "00000000";
IM(4194388) <= "10110011";
IM(4194389) <= "00000110";
IM(4194390) <= "00000101";
IM(4194391) <= "00000000";
IM(4194392) <= "11101111";
IM(4194393) <= "11110000";
IM(4194394) <= "01011111";
IM(4194395) <= "11111100";
IM(4194396) <= "00010011";
IM(4194397) <= "00000000";
IM(4194398) <= "00000000";
IM(4194399) <= "00000000";
IM(4194400) <= "00010011";
IM(4194401) <= "00000000";
IM(4194402) <= "00000000";
IM(4194403) <= "00000000";
IM(4194404) <= "00010011";
IM(4194405) <= "00000000";
IM(4194406) <= "00000000";
IM(4194407) <= "00000000";
IM(4194408) <= "00100011";
IM(4194409) <= "10100000";
IM(4194410) <= "11010010";
IM(4194411) <= "00000000";
IM(4194412) <= "11101111";
IM(4194413) <= "00000000";
IM(4194414) <= "00000000";
IM(4194415) <= "00000000";
IM(4194416) <= "00010011";
IM(4194417) <= "00000000";
IM(4194418) <= "00000000";
IM(4194419) <= "00000000";
IM(4194420) <= "00010011";
IM(4194421) <= "00000000";
IM(4194422) <= "00000000";
IM(4194423) <= "00000000";
IM(4194424) <= "00010011";
IM(4194425) <= "00000000";
IM(4194426) <= "00000000";
IM(4194427) <= "00000000";


--IM(4194504) <= "00010011";
--IM(4194505) <= "00000000";
--IM(4194506) <= "00000000";
--IM(4194507) <= "00000000";

--IM(4194508) <= "00010011";
--IM(4194509) <= "00000000";
--IM(4194510) <= "00000000";
--IM(4194511) <= "00000000";

PROCESS(CLK)
VARIABLE DATA_OUT_s: STD_LOGIC_VECTOR(31 DOWNTO 0); -- USING A VARIABLE TO AVOID TIMING ISSUES
BEGIN


	IF(CLK'EVENT AND CLK = '1') THEN
		IF (MEM_READ = '1') THEN
			IF (TO_INTEGER(UNSIGNED(ADDR))>4194428 OR TO_INTEGER(UNSIGNED(ADDR))<4194300) THEN
				DATA_OUT_s := (OTHERS =>'0');

			ELSE
				DATA_OUT_s := IM(TO_INTEGER(UNSIGNED(ADDR)+3)) & IM(TO_INTEGER(UNSIGNED(ADDR)+2)) & IM(TO_INTEGER(UNSIGNED(ADDR)+1))
								& IM(TO_INTEGER(UNSIGNED(ADDR))); --LSBytefirst
			END IF;

			DATA_OUT <= DATA_OUT_s;
		END IF;

	END IF;

END PROCESS;

END structure;
